module part2 (SW, HEX1, HEX0);
    input [3:0] SW;
    output [0:6] HEX1, HEX0;
endmodule