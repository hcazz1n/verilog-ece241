module part1 (SW, LEDR, HEX1, HEX0);
    input [7:0] SW;
    output [7:0] LEDR;
    output [6:0] HEX1, HEX0;
endmodule