module part4 (SW, LEDR, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0);
    input [8:0] SW;
    output [9:0] LEDR;
    output [6:0] HEX5, HEX4, HEX3, HEX2, HEX1, HEX0;
endmodule